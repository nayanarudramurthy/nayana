module gui();

endmodule
