module radhika()

endmodule
