module nayana()

endmodule
