module radhika()

endmodule :
